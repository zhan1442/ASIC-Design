/home/ecegrid/a/mg112/ece337/Lab2/source/tb_adder_nbit.sv