/home/ecegrid/a/mg112/ece337/Lab2/source/adder_nbit.sv